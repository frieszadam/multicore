`ifndef CORE_VH
`define CORE_VH

// Defined in the OpenHW-OBI specification for atop signal
`define ATOP_LR 5'h2
`define ATOP_SC 5'h3


`endif
